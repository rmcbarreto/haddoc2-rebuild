library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.math_real.all;
library work;
use work.cnn_types.all;

entity DotProduct is
  generic(
    BITWIDTH       : integer; -- 8
    SUM_WIDTH        : integer; -- 3*8 -> 3*bitwidth
    DOT_PRODUCT_SIZE : integer; -- KERNEL_SIZE*KERNEL_SIZE
    KERNEL_VALUE     : pixel_array; -- gets the values from params
    BIAS_VALUE       : std_logic_vector
    );
  port(
    clk      : in  std_logic;
    reset_n  : in  std_logic;
    enable   : in  std_logic;
    in_data  : in  pixel_array (0 to DOT_PRODUCT_SIZE - 1);
    in_dv    : in  std_logic;
    out_data : out std_logic_vector (SUM_WIDTH-1 downto 0);
    out_dv   : out std_logic
	 --out_aux_data   : out std_logic_vector(7 downto 0);
	 --aux_dv	 : out std_logic
    );
end DotProduct;

architecture rtl of DotProduct is
  --------------------------------------------------------------
  ---- Implementation with the multiplier and adder components
  --------------------------------------------------------------
  component MCM
     generic (
       BITWIDTH       : integer;
       DOT_PRODUCT_SIZE : integer;
       KERNEL_VALUE     : pixel_array
       );
     port (
       clk       : in  std_logic;
       reset_n   : in  std_logic;
       enable    : in  std_logic;
       in_data   : in  pixel_array (0 to DOT_PRODUCT_SIZE - 1);
       in_dv  	  : in  std_logic;
       out_data  : out prod_array (0 to DOT_PRODUCT_SIZE - 1); -- prod_array -> 2*GENERAL_BITWIDTH = 2*8
       out_dv 	  : out std_logic
       );
  end component MCM;
  --
  component MOA
     generic (
       BITWIDTH   : integer;
       SUM_WIDTH    : integer;
       NUM_OPERANDS : integer;
       BIAS_VALUE   : std_logic_vector
       );
     port (
       clk       : in  std_logic;
       reset_n   : in  std_logic;
       enable    : in  std_logic;
       in_data   : in  prod_array (0 to NUM_OPERANDS - 1); -- prod_array -> 2*GENERAL_BITWIDTH = 2*8
       in_dv  	  : in  std_logic;
       out_data  : out std_logic_vector (SUM_WIDTH-1 downto 0);
       out_dv	  : out std_logic
       );
  end component MOA;
  --
  signal p_prod_data  : prod_array (0 to DOT_PRODUCT_SIZE - 1);
  signal p_prod_valid : std_logic;
  
  --signal aux_aux : std_logic_vector(15 downto 0);
  
   begin
	
	--aux_dv <= p_prod_valid;
	
	--aux_aux <= To_StdLogicVector(out_data(4));
	--out_aux_data <= aux_aux(7 downto 0);
	--out_aux_data <= p_prod_data(8)(7 downto 0);
	--out_aux_data <= out_data(7 downto 0);
	
   MCM_i : MCM
     generic map (
       BITWIDTH       => BITWIDTH,
       DOT_PRODUCT_SIZE => DOT_PRODUCT_SIZE,
       KERNEL_VALUE     => KERNEL_VALUE
       )
     port map (
       clk       => clk,
       reset_n   => reset_n,
       enable    => enable,
       in_data   => in_data,
       in_dv	  => in_dv,
       out_data  => p_prod_data,
       out_dv	  => p_prod_valid
		 --out_dv	  => out_dv
       );
		 
   MOA_i : MOA
     generic map (
       BITWIDTH   => BITWIDTH,
       SUM_WIDTH    => SUM_WIDTH,
       NUM_OPERANDS => DOT_PRODUCT_SIZE,
       BIAS_VALUE   => BIAS_VALUE
       )
     port map (
       clk       => clk,
       reset_n   => reset_n,
       enable    => enable,
       in_data   => p_prod_data,
       in_dv	  => p_prod_valid,
       out_data  => out_data,
		 out_dv	  => out_dv
       );
   

  --------------------------------------------------------------
  ---- Direct Implementation as a Pipelined MAC
  --------------------------------------------------------------
--  signal pip_acc : sum_array (0 to DOT_PRODUCT_SIZE - 1) := (others => (others => '0'));
--  begin
--    process(clk)
--    begin
--      if (reset_n = '0') then
--        pip_acc <= (others => (others => '0'));
--        out_dv  <= '0';
--        out_fv  <= '0';
--
--      elsif(rising_edge(clk)) then
--        if (enable = '1') then
--          if (in_dv = '1' and in_fv = '1') then
--            pip_acc(0)(2*BITWIDTH-1 downto 0) <= in_data(0) *  KERNEL_VALUE(0);
--            acc_loop : for i in 1 to DOT_PRODUCT_SIZE-1 loop
--              pip_acc(i) <= pip_acc(i-1) + (in_data(i) * KERNEL_VALUE(i));
--            end loop acc_loop;
--          end if;
--          out_dv <= in_dv;
--          out_fv <= in_fv;
--        end if;
--      end if;
--    end process;
--    out_data <= pip_acc(DOT_PRODUCT_SIZE-1) + BIAS_VALUE;
end architecture;
