------------------------------------------------------------------------------
-- Title      : convElement
-- Project    : Haddoc2
------------------------------------------------------------------------------
-- File       : convElement.vhd
-- Author     : K. Abdelouahab
-- Company    : Institut Pascal
-- Last update: 2018-08-23
------------------------------------------------------------------------------
-- Description: A fully pipelined implementation of CNN layers that is able to process
--              one pixel/clock cycle. Each actors of a CNN graph are directly mapped
--              on the hardware following the principals of DHM and DataFlow processing
--                            ______
--                          |       |
--                          |       |-- output_streams-->
--        input_streams---->| conv  |-- output_streams-->
--        input_streams---->| Layer |-- output_streams-->
--        input_streams---->|       |-- output_streams-->
--        input_streams---->|       |-- output_streams-->
--                          |       |-- output_streams-->
--                           ______
-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.math_real.all;
library work;
use work.cnn_types.all;
--==================================================================
-- Added by, Ricardo Barreto
use ieee.numeric_std.all;
--==================================================================


entity ConvLayer is
  generic(
    BITWIDTH   : integer;
    IMAGE_WIDTH  : integer;
    SUM_WIDTH    : integer;
    KERNEL_SIZE  : integer;
    NB_IN_FLOWS  : integer;
    NB_OUT_FLOWS : integer;
    KERNEL_VALUE : pixel_matrix;
    BIAS_VALUE   : pixel_array
	 
--    BITWIDTH   : integer := 8;
--    SUM_WIDTH    : integer := 3 * 8; -- 8 is the general bit width
--	 IMAGE_WIDTH  : integer := 28;
--    KERNEL_SIZE  : integer := 3;
--	 --KERNEL_SIZE  : integer := 3;
--    NB_IN_FLOWS  : integer := 1; -- number of inputs (if greyscale 1 input, if colormode RGB 3 inputs)
--    NB_OUT_FLOWS : integer := 1; -- number of convolutions
--    --KERNEL_VALUE : pixel_matrix	(0 to NB_OUT_FLOWS - 1 ,  0 to NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE - 1) :=
--	 --KERNEL_VALUE : pixel_matrix	(0 to 1,  0 to 24) :=
-- --( ("00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001"),
--	--("00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001")
--	--);
--	KERNEL_VALUE : pixel_matrix	(0 to 1,  0 to 8) :=
-- ( ("00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001"),
--	("00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001")
--	);
--    --BIAS_VALUE   : pixel_array	(0 to NB_OUT_FLOWS - 1 ) := ("00000001")
--	 BIAS_VALUE   : pixel_array	(0 to 1 ) := ("00000001", "00000001")
    );

  port(
    clk      : in  std_logic;
    reset_n  : in  std_logic;
    enable   : in  std_logic;
    in_data  : in  pixel_array(0 to NB_IN_FLOWS - 1);
    in_dv    : in  std_logic;
    out_data : out pixel_array(0 to NB_OUT_FLOWS - 1);
    out_dv   : out std_logic
	 --aux_out	 : out std_logic_vector(15 downto 0); -- used for things like counters
	 --aux_out_dv : out std_logic; -- tensorExtractor
	 --aux_out_fv : out std_logic;
	 --aux_out_data_test : out pixel_array(0 to (KERNEL_SIZE*KERNEL_SIZE-1)); -- tensorExtrator
	 --out_aux_data   : out std_logic_vector(7 downto 0) -- dotProduct
    );
end entity;

architecture STRUCTURAL of ConvLayer is
  --------------------------------------------------------------------------------
  -- COMPONENTS
  --------------------------------------------------------------------------------
  component TensorExtractor
    generic (
      BITWIDTH  : integer;
      IMAGE_WIDTH : integer;
      KERNEL_SIZE : integer;
      NB_IN_FLOWS : integer
      );
    port (
      clk      : in  std_logic;
      reset_n  : in  std_logic;
      enable   : in  std_logic;
      in_data  : in  pixel_array (0 to NB_IN_FLOWS - 1);
      in_dv    : in  std_logic;
      out_data : out pixel_array (0 to NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE- 1); -- 0 to 1*3*3 -1  = 9 elements
      out_dv   : out std_logic
      );
  end component TensorExtractor;

  component DotProduct
    generic (
      BITWIDTH       : integer;
      SUM_WIDTH        : integer;
      DOT_PRODUCT_SIZE : integer;
      KERNEL_VALUE     : pixel_array;
      BIAS_VALUE       : std_logic_vector
      );
    port (
      clk      : in  std_logic;
      reset_n  : in  std_logic;
      enable   : in  std_logic;
      in_data  : in  pixel_array (0 to DOT_PRODUCT_SIZE - 1);
      in_dv    : in  std_logic;
      out_data : out std_logic_vector (SUM_WIDTH-1 downto 0);
      out_dv   : out std_logic
		--out_aux_data   : out std_logic_vector(7 downto 0)
      );
  end component DotProduct;


  component TanhLayer
    generic (
      BITWIDTH : integer;
      SUM_WIDTH  : integer
      );
    port (
      in_data  : in  std_logic_vector (SUM_WIDTH-1 downto 0);
      out_data : out std_logic_vector (BITWIDTH-1 downto 0)
      );
  end component TanhLayer;
  
  
------------------------------------------------------------------------------------------
  signal neighborhood_data : pixel_array (0 to NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE- 1); -- 0 to 1*3*3 -1  = 9 elements
  signal neighborhood_dv   : std_logic;
  signal dp_data           : sum_array (0 to NB_OUT_FLOWS-1);
  signal dp_dv             : std_logic;
-----------------------------------------------------------------------------------------

begin

--aux_out_data_test <= neighborhood_data; -- tensorExtrator

--aux_out_dv <= neighborhood_dv; -- tensorExtrator


  TensorExtractor_i : TensorExtractor
    generic map (
      BITWIDTH  => BITWIDTH,
      IMAGE_WIDTH => IMAGE_WIDTH,
      KERNEL_SIZE => KERNEL_SIZE,
      NB_IN_FLOWS => NB_IN_FLOWS
      )
    port map (
      clk      => clk,
      reset_n  => reset_n,
      enable   => enable,
      in_data  => in_data,
      in_dv    => in_dv,
      out_data => neighborhood_data, -- output array of 8 bits with size of 9 elements
      out_dv   => neighborhood_dv
		--out_dv   => out_dv
      );

		
  DotProduct_loop : for n in 0 to NB_OUT_FLOWS- 1 generate
  
  --==================================================================
  -- Added by Ricardo Barreto
	first_Dotproduct : if n = 0 generate
    DotProduct_i : DotProduct
      generic map (
        BITWIDTH       	 => BITWIDTH,
        SUM_WIDTH        => SUM_WIDTH, -- 3*8 -> 3*bitwidth
        DOT_PRODUCT_SIZE => NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,
        BIAS_VALUE       => BIAS_VALUE(n),
        KERNEL_VALUE     => extractRow(n,
                                   NB_OUT_FLOWS,  -- N
                                   NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,  -- CJK
                                   KERNEL_VALUE)  --Theta(n)
        )
      port map (
        clk      => clk,
        reset_n  => reset_n,
        enable   => enable,
        in_data  => neighborhood_data,
        in_dv    => neighborhood_dv,
        out_data => dp_data(n),
        out_dv   => out_dv
		  --out_aux_data   => out_aux_data
        );

    -- Dummy Activation
    TanhLayer_i : TanhLayer
      generic map (
        BITWIDTH => BITWIDTH,
        SUM_WIDTH  => SUM_WIDTH
        )
      port map (
        in_data  => dp_data(n),
        out_data => out_data(n)
        );
		  
	end generate first_Dotproduct;
	
	other_DotProduct : if n > 0 generate
		DotProduct_i : DotProduct
      generic map (
        BITWIDTH       => BITWIDTH,
        SUM_WIDTH        => SUM_WIDTH,
        DOT_PRODUCT_SIZE => NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,
        BIAS_VALUE       => BIAS_VALUE(n),
        KERNEL_VALUE     => extractRow(n,
                                   NB_OUT_FLOWS,  -- N
                                   NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,  -- CJK
                                   KERNEL_VALUE)  --Theta(n)
        )
      port map (
        clk      => clk,
        reset_n  => reset_n,
        enable   => enable,
        in_data  => neighborhood_data,
        in_dv    => neighborhood_dv,
        out_data => dp_data(n),
		  out_dv   => open
		  --out_aux_data   => open
        );

    -- Dummy Activation
    TanhLayer_i : TanhLayer
      generic map (
        BITWIDTH => BITWIDTH,
        SUM_WIDTH  => SUM_WIDTH
        )
      port map (
        in_data  => dp_data(n),
        out_data => out_data(n)
        );
	end generate other_DotProduct;
	
--==================================================================
	
	
	--==================================================================
	-- ORIGINAL
--	DotProduct_i : DotProduct
--      generic map (
--        BITWIDTH       => BITWIDTH,
--        SUM_WIDTH        => SUM_WIDTH,
--        DOT_PRODUCT_SIZE => NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,
--        BIAS_VALUE       => BIAS_VALUE(n),
--        KERNEL_VALUE     => extractRow(n,
--                                   NB_OUT_FLOWS,  -- N
--                                   NB_IN_FLOWS * KERNEL_SIZE * KERNEL_SIZE,  -- CJK
--                                   KERNEL_VALUE)  --Theta(n)
--        )
--      port map (
--        clk      => clk,
--        reset_n  => reset_n,
--        enable   => enable,
--        in_data  => neighborhood_data,
--        in_dv    => neighborhood_dv,
--        in_fv    => neighborhood_fv,
--        out_data => dp_data(n),
--		  out_dv   => open,
--        out_fv   => open
--        );
--
--    -- Dummy Activation
--    TanhLayer_i : TanhLayer
--      generic map (
--        BITWIDTH => BITWIDTH,
--        SUM_WIDTH  => SUM_WIDTH
--        )
--      port map (
--        in_data  => dp_data(n),
--        out_data => out_data(n)
--        );
--    out_dv <= in_dv;
--    out_fv <= in_fv;
	 --==================================================================
  end generate;



end architecture;
